`default_nettype none

module pixel_ram_block(
    input wire i_clk,
    // Write interface
    input wire [7:0] i_w_addr,
    input wire [15:0] i_w_data,
    input wire i_w_enable,
    // Read interface
    input wire [7:0] i_r_addr,
    output reg [15:0] o_r_data,
    input wire i_r_enable
);

reg [15:0] data[256];
integer i;
initial begin
    for (i = 0; i < 256; i++)
        data[i] = 16'h80;
end

always @(posedge i_clk)
    if (i_r_enable)
        o_r_data <= data[i_r_addr];

always @(posedge i_clk)
    if (i_w_enable)
        data[i_w_addr] <= i_w_data;

/*

SB_RAM40_4K #(
    .READ_MODE(0), // 256x16
    .WRITE_MODE(0), // 256x16
    .INIT_0(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_1(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_2(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_3(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_4(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_5(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_6(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_7(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_8(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_9(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_A(256'H00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000)
) ram40_upper (
    .WADDR(i_w_addr),
    .RADDR(i_r_addr),
    .MASK(16'b0), // 0 = write, 1 = don't
    .WDATA(i_w_data),
    .RDATA(o_r_data),
    .WE(i_w_enable),
    .WCLKE(1'b1),
    .WCLK(i_clk),
    .RE(i_r_enable),
    .RCLKE(1'b1),
    .RCLK(i_clk)
);

*/
    /*
    .INIT_0(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
    .INIT_1(256'h11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111),
    .INIT_2(256'h22222222_22222222_22222222_22222222_22222222_22222222_22222222_22222222),
    .INIT_3(256'h33333333_33333333_33333333_33333333_33333333_33333333_33333333_33333333),
    .INIT_4(256'h44444444_44444444_44444444_44444444_44444444_44444444_44444444_44444444),
    .INIT_5(256'h55555555_55555555_55555555_55555555_55555555_55555555_55555555_55555555),
    .INIT_6(256'h66666666_66666666_66666666_66666666_66666666_66666666_66666666_66666666),
    .INIT_7(256'h77777777_77777777_77777777_77777777_77777777_77777777_77777777_77777777),
    .INIT_8(256'h88888888_88888888_88888888_88888888_88888888_88888888_88888888_88888888),
    .INIT_9(256'h99999999_99999999_99999999_99999999_99999999_99999999_99999999_99999999),
    .INIT_A(256'HAAAAAAAA_AAAAAAAA_AAAAAAAA_AAAAAAAA_AAAAAAAA_AAAAAAAA_AAAAAAAA_AAAAAAAA),
    .INIT_B(256'hBBBBBBBB_BBBBBBBB_BBBBBBBB_BBBBBBBB_BBBBBBBB_BBBBBBBB_BBBBBBBB_BBBBBBBB),
    .INIT_C(256'hCCCCCCCC_CCCCCCCC_CCCCCCCC_CCCCCCCC_CCCCCCCC_CCCCCCCC_CCCCCCCC_CCCCCCCC),
    .INIT_D(256'hDDDDDDDD_DDDDDDDD_DDDDDDDD_DDDDDDDD_DDDDDDDD_DDDDDDDD_DDDDDDDD_DDDDDDDD),
    .INIT_E(256'hEEEEEEEE_EEEEEEEE_EEEEEEEE_EEEEEEEE_EEEEEEEE_EEEEEEEE_EEEEEEEE_EEEEEEEE),
    .INIT_F(256'hFFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF)
    */

endmodule
